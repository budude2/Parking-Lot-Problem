`timescale 1ns / 1ps

module lotTracker(

    );
endmodule