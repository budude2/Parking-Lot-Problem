`timescale 1ns / 1ps

module carCounter(

    );
endmodule
